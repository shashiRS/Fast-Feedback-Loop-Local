MIIJiwYJKwYBBAGCN1gDoIIJfDCCCXgGCisGAQQBgjdYAwGgggloMIIJZAIDAgAB
AgJmAQIBQAQIz11sn9FkpKYEEF1edKUjMd9LiSEsR4eRWBAEggk4p1Vaf4U1jprW
AIxjbn4Q1lg9EUmSEy1dcoSiRvyP16KpHrsk/dBvHwGm/Xwdg+tdJdKfEB/Cdrkt
PxBa3BEt9Ow+SyLyU++GclN5S5LhvGc2nHvhGX6or6Zspyjq2y/7lAPxlMnvUXoY
tTtl9BwBNDMt9T4yNRqP2RMgpaGqsUJdg75QL9gGjCXt+FZm1li90hD6QXOg3xFK
DI18Y1johoRYinnOJsJApZDw6nkmnkgBFEFofiALxyF3M96ckPB9wdLRER6tTv7l
9EklUHdszbQcU79upkJt8WeQFmbX4tQSPacwMX0abh661KRV/ECxz2AtyMpsXkVp
lQCjCddInUoShKEb7qVcZuTcaBNJS5PoUj3tWXbaEwBadK4peOkJVuGhfhhUM9gA
7CPikt4a731LJ0zDfJlztLcLtq57+lOYdMW9x/g1v9IZ1X5hLqc/inI1nQNifxqn
R6r2ZskvQgZwGXxXbQR7tImISUGfiTuaydUNR77m6f45jLLoC5rWjvZawyWdP44X
KnxINxOynOq7tinHudw+0EDrDS8/IPYYknqupZlJ0b56Ov8Q/4A7C0UmLeloTFdk
SRI1vzWrwVSD+pXM5wTTWmpMcQtoD5kSXC3mYRGCRIk3ZXs4dQ2nmXN9fDQJQMbG
aZfL0SRNe3mDKfl8MQ+G0n5j+rVWaOK8ZJwqYIblEZHBiM0pJZELCclRapGQ0pX3
YhH71vImM+f8dPLZf7WK6UF6eL/M5XuEGce9K2lE9UIUrR72aNpYWV/05TCug+mi
qz8GSpoCTgjwQHy06Z1nYT++qDzauAeOerYAdZH11JlSNEgA1qqHbxPjq53FRQUH
1BSRigVyYV0qlAMs/X1zNo0as7cwX0L/165vgBb3dBw6b0aE7M3M7FYt99b9NPMM
8lx/AaZINn0founhcJ9r1RV3IrrT6ugIFS04wfN8aCEAiOpIiSmu/63SwAn6U+QK
KRJvYiXhLbYZRszYnVugxokLEYCzu0CvIGCTcgYtxOYdKvl743TQfJ4AAhIVPy5p
F60fOnhZD0eORz+PBiM2q9CH+SQVB+FYMb8mvV7rOIxAAEdbba4x4b79wJMPMrN2
QT4gMYiWJYTEcCOupwcFJcKJlTLgb2lIpnUllHDx1M8hrePRBjtyVPJv8w+JqG9F
/b1VAiT8fQEyBlaq118Z3oNosLwgEhcDhiC/wWhvVGcbgtq66ametc2Xv4+8CVdb
hml7wt5SUkLXDP6B5WC9UJwYt3+6bA0nOoFF23X2a5ViVQh3yBlLgLZTppyHyBub
cGosQC8T3HuV8Os9Lv8vCNpavEaGGvejEBuYi9sRu5vNem2EtdrCbYYS1U+EI0/j
SccXLXUq9HI4d3TAYZxBZKPGJqQCkdfYQq4fpKs3OjV6vmndKefZfgxbE5+1gFGQ
kkgjABMjxOLFbdx2P4u0480fffOPF2XapE3kl6ZnSIC/4DETimvCnt6d0pUiM6fB
hIxorGP1iXSQzCH5PcDo5NkBmI9MSvBiuk01LN5cHfTGfZcMdBNls683n+qhm5x6
SJCWYTd7T5Fcjm/3qZMNtklNw7eQgvlQfcu7cvycfyDQ8lTNzT8Cq6huj97OH1kb
iPm78Koz10TxezA++zP4zLjrUEG/UC11e54+LtJv0zKmlfy3OAqndvYwtyR4RjhQ
kBFNJGCwjlGXN1m/1GYfe7o7o/QATrjB+MJ62wOora9isSPY4h560q15kHU8FoeP
KhSLbznijjnFLuAu1OUjgQnTqwEgiAUDM+seZS96gQMgsePaBAOhmTqTEesSVWwn
Cfx5slzi3Jxm0b+P4EvenH53WvCAowHsYrnyDHdsEM++GslwRVqVGMltfUAUCMyi
tEZpHMiPC4sSEv+EOmVLRc1Y5ts03qCdbuiRgA+XKAJ+8NGeg5DNJwncUZlsOxQd
/HrBcAsHN+VKfmF2BZeiQuZYFP0wnZnqwImHaSvcB9QWBNFT1/qyzZcS6yNYvUGw
zlW7SuA1II5Zi6yZ6W+HCa7tdW6ifGWTiwds4TxxtABO7SCDYLMLkm+Z6l/4GpOk
PrZGK54msOLgj/a8iVYYNP7kLAFsEcF53gRSddQ7Fj9lrDktg8GzZWIXOGIjx7ae
PKMxYKOGIGfc0bLMH5t4+j0+0ZitxeCeuvK2p0fztqAD432ZFyg5oQXvScWXBtLn
RxfwEjdPEVHY99eFZi41qdpRuQ5xB80r6e2/2O4MMQD4fkm1zfPhybNkELFy51in
krlP0MpXVC+zpIfePTzUkMgOvPQg+S9Lrrryx3SjZT9uDABoS+1v4pmetSJZCmXR
AddO3LyNb6FGMrpC9MQBYtItptFcnoOQHg0zw0yWu8z6JR0nAk5wxZPICfND1KKe
bffOsKOHwVqgbyH9uC61m7nUHcsPoUbykwgVWdA8zyPcAUJgfcl36w7N5TImA0Ok
K7gEjgNN9/iQXmcJPaKUQkwV7hBDj2AVOt0rNU6f926DFcPe3IB3w7Vg+9FO6Uj9
YeHNjDmipjZmbk3wURZYEDz4HtKNEzXpqzUSvA2//b9IMFQgSiGqz++6SDjgQP3V
++6/Y3sSyUCX4Ub93K4rwvcfh74ghccctrlFt5ul/Z2NWOS0rySYA86ou02HlONj
NSvjw74EVqzksQZMcwyXP6iuHy+tYOpeGAY6uuPbBz9oulwL6rZAj1OWOWy6GeNz
cLfLxv6SKyULJz4KsBJUgyduQAVkglXz7hqoItFAqUy3tDLVlV1jvpZcbEm6bqWT
QTsAe7KB0i/prwMeDdSvSfQnq4eW7g0EoGWq0qvLChOEsabWyfItJekG11PcHDw9
e6/tVSMR2bA+QWtU28Bs4iruTB1tSqvWhLSNrM8cax/RXWPvHV6+tERw0aKqGasW
1f6B13xPyuCv6jyW1MAkHJrE5deUbflesuXPnTzCcuGpijiKGUvMlS3p2EVd3QKm
PN+78tjuhKMCLcHmEzIPE1clwKlvYWZgbUPj0xnkFJ21/+2L1IhIEI1TO/dxfalp
x2VqK+3diSwSGadQ+/EhM0EnD+ftSrRP/0TYrNcuGFpbdI5YSUFpuQPSEvoPK5JL
5ErIwYdBC+pJQC+2Q4hdWSsM9AvVLbLkhVgC5IqynRCD0QzIn5kTQtn/JiI+UAU=
MIIJiwYJKwYBBAGCN1gDoIIJfDCCCXgGCisGAQQBgjdYAwGgggloMIIJZAIDAgAB
AgJmAQIBQAQIoZWClcMxDIwEELQh03EgJZ8f4+XLdt0ho7oEggk4W7meHWnuGpdm
b4hTjPDXbvQ9oZcPTCPxBccMcFqApX3YL0Wq33k5Z+mfQf11/ZXHDLGMAYVjXCKr
bXknKsTczlWr0dpAwVlAaeUnIn6Xkg+8RfKKjT9xYx20Gi0o2O5ug0mmZr3+tloK
zvoD8Fc18xdQg6BFAjc0OvrldqNh1nF4/KZNDMB//Z0sgzt+uKEZRSaPYXw+qvud
qcTvG1kzea9+S9KVEdItpcAoUl8Njr6ccL27AERoC98/IEr0dg7cEa/28qPY+zzG
upPpA+k0AFy6AKH6h6MbQKg2Ew3yEW+5a2y0nUJUVasTzhjzwVxXITcwn/97d2QA
O5pKtxcDz1bwZXwkcj1GhYE+0LWLlR7yyHtSCo4CJX5tA5p5ObhAbkZhA6uvdcDa
hkzGvC2BgObnDS/AcUjASV8FN1HZBLtzGfxshzF4KZN0AF+n04uIEUbVLCuJ/lnW
q0V3XKUqYMJXBtAzxlcu76KcjDv2FBTRj22kaAnADwvOhmSrDGHj+LoUIhO/fiWH
fsgokNo7JlOSyodsRvcbmqFiEih6avSUm2INbQofUuA0jKmoFdtQ7TJ4EOWhx52Z
PGgdeJxKve83yOQQsRHwOXV3plMZuSVYWNuxTODC2xJISKZYteyu9ct4OX+pmjw4
CUChqem2MaYGCaPolxR0IaVvCR1tD2llfpbuSeuS3TFTajb7OMJm+2jqJtGpLbsO
K6ZmC6Y7ooNmmJphwLmd3V2Y86oQi3fJOCgmS8kKbCs9UXNH4+u8z1sILcOdlXqG
2xeRHt902iRIWx9QhIkhFd06CsuuBdZnDqj7Mu/pkh7KmHOpM12X//i+83k1cFRb
oaqjney8XbzoqqvjVpu10IrwvIB17jt/Pw4B5H5thLgJBcBMSRur3qK5V8I7adM2
81Z3Nu+1tm0LotOMtGEEi/hCvwgOiOWUtqsC1anqkyISm6lCMEMSctEa50rGaw/8
lMy1o8KUYOpWLKB2RTZ/mR9SlAH7HWotX9Fuk8HGwZE3lyyADayh2T39BNl2yDk/
JUmNh3HsXi6PPogKdLbyX0TBImFxCEfOLGbL62CZ1PKXsgzbviIrc6GJ08wEDS0j
KdGIV3Pfovvn30uWfh/vSOypDZx8+wI105F+BBJEg+inXjjSI4qZz97hmco8m1nP
nOmjolJhNsjhea/46W5BfztUmXvJyjbVNiYTW5U27j9rylgD6myMQBptEJ79dPio
haMc7ifTUiua/UW91RGEIjYb0g3HWVsGQbVhZ3Y1CDPBA6FBE6PVOjTBEyZ11Q89
lX2cB2CSSMQXXFLVQc8MYA8IjTD3ekoed7hH1205LSwvkYN+ycJKPRtzHDDU6RZu
mNXghbW2Ez0lLcu8B6Ei9Ew/Jyog2UcFxyCiY5abvc/qM7l5TUCBsG3R7MzQ+t5C
zTdZiAEuMNyskZC73qAvtWhzyaVKd8bWV9EsFUOylDYL/yVH8sw99NWjtQnK7mmN
RPOLR8r7YT8JOKmz3GOmQYVDOqR9Gv4mUS4Wf78h4TkX5ozk0J+qP3ioSkbp4LE0
SrG58xz2YEN7705fgK56LQ1RnibaSU2S06Kzz7ew9rrUkJropeLjz8znfjyQHzYd
O1jKPm/1yC+fZWpfI4BCDJWh1gtqTt8GIq6N4PHteP+4NAeX1PJh1hnILK+WPmyW
jNHLz16OW+XBCaEDOiC8m+ukzmzd2BfzNDQP3OJrPlUItJ1OGpZfZl8lockm/Zrb
IICo+qG1ezGeS6UDBSIFz5xyk5ksQw8MlhsdDS/XEP/GapomAUvmi3FQ6moF3lPi
5dKo7fwUEnurPtCPFolpN24pibC550F+GzuaLv4VNB5FT6ZmqnJFvwGelz7vIGVt
q3Hwk0a6xjJoMhvEaWgPO7EHwCqKPr6pJKXX4Fxznx9LncxqqFLHuHuz/BcxGIIj
8pWXRcfXYHY9W5J6Azo9I5JA4K/coKSlRsTwJ88Vz1xRylFRoFf/hF9XNyBAAho8
rN4emuCq5jFwHXvtoPXO/DODKusJm5GXev4yO8v5YMZoC0Xz00YtMpRni0lZZr09
pJCTsZCD1tSM3VeVfJ0hOg0VFssx6RFjq5QIdT6rosMEvbNx6G6MswPCmnCxjk+m
z+u1S1fOvGfAohb20jWt5Vr3+/M+1kbKJqOFNFVsOEvXdJN4eba6um6nsAYchQJu
eY6LmBtVvIMq5pHI1EIucOf3CiLOF/c4tCw5ze33b0EHwYD5LSkWFOEiPeyMO6sZ
ULlc1UcAr6NXdMhIgSU2diYiqRnKCMJPkwhwcfEjNGWyQefdkPLKYuLpVjDeIWf/
bdMpLFhm70BFMo/HMupbhrmchV8p5EULC9sWOkMqGYREDUQnfGrYBFlMeO9gfiGq
tN1266RBd2ES4/AyX8+Ftr811LrTkSzSTx6LQDKIewQLD3OszNpmZTgepeCAfbKK
mIuN47re4VcZqVgu9z0ixy/NqEo6ljIH5j5RtjVmAGgmqbX7+iNik568ydedCIIa
UPiKoGP3w1hoYHONGNM1RniVPOkdk64TpfqhpQ02EftsGBokKP/B8PA2d2c8THVn
AS5wKpOFsJN7Rb133w3pi8OZq08Bkz8f71xefQzifiI33Rk1IZEyC9UBOgCS7bVj
+k3Rs527G0VSlZZ/Lf+czp/4jpPEL/LF8JYLEIH/DST9q2zdK4uxZHTh39UEr5QL
n6upIfjsmajbqEqGEKaaWGu54/0KTBFOUCB00ymSoBWgsnYPK8BJLKH4bVn71wX2
apzUZUx5KPuTBlDFPf6SFJIc3Xgm4TfbhJy4qkqV2ljQcDctFyLhOIllFhqzb+Wx
o/yQMVDqDnSsxVipatebOzvuz7caIjBa4dBknOWxSS+m6hW8JHkWZYngQkFISwWd
Uno6ApNIb2Tl1y1/m7L+9ZhxM0O6BQeA4MRnmRQ4XF4BwxD6TYi9OhODvbpY3yiY
3JvcZz7Y0KMpS6a+XmVxq1g40Gu0rvCrouS5IzLDDPcDBIKRfzTrSqbJg/lFSGlP
BVADQLmPLLKmZwPZ46S32D++ycDc7GMOOK0II+XT1SF3wsVeLQR9gwv7B1MdSafK
ge5UUhds8Xs3ZJBsUnGzkWvpzXOeZARbCCMmQt+1WCpNDtqpiYhPIIBb8I6MLLU=

MIIIowYJKwYBBAGCN1gDoIIIlDCCCJAGCisGAQQBgjdYAwGgggiAMIIIfAIDAgAB
AgJmAQIBQAQI2L0cmJRdvQQEEKlAWijma7HQvNr8WNXhDJgEgghQ3p6YylRtavaH
XShFs+ysdZt+LE86Px0ippjZtwyxEzeUDECNupNsxlxzt4/vmaYuP81EUGjKvV3Q
HmLvu0xCByHX4P2EBwKqy5PeQChGiyVkH4SVALxusvW8jgNQQdkBrccCc5O4jqgD
o57wP36F+Si+rTSexixNb9wlpXqBax2qC4bl54EwOn/QbTNE4h79MVMihAdHY/5b
xBbINpIfL7/LlO/F5taRfxOWYeyk8AfuWUXBGpB+2YnkYZIWU/Dk5NJAxE0Pnb4U
S7644DBFWUWbjEfu9jxZsTEVBim6fv/dJ3lSyTE3Wsj7IL2RQuDmR30ZgzQVrulu
N0wRm8wSC8aoclaFPnZh7atCiYJCC2LjzXxuUbs+DJvg1eMu0PnahE4NumwFN0Rt
0DC9nq8JcJuuneOLisbe90Blm15SZdXH9Yqz/Q5Wvd6wq1wiA67V7Uri1hASlFrv
0WpB1k4/o9mpiFT173d8CrzWZNivsaxPgKUnDX+LA2Txb3QMnVhB7LpOCl0Qnwwt
O1+NhPoLUE2v3J8s0UD7puKfXCgXjiSb7xvFPbdBfmgKvaHxrb35NJK7GGq8VXJG
Sq++pV/kBoNtWhO1zwSJ9cV0N5umsnSlbYaduQmmZVFCHXnhpOxi3uZ2PS+3TmSR
V07r5zPV47zE+8fMeFW5PY6Qtv5q6ce2uEYFWkoy4gHmCPCEDxznYEMPsYeozOrS
iXMxfteR64oAz9oTn4FRQlgnsMfBheGndi3jHfgx0VT3HCw9u9UZ0kugwXZmsmKM
JYfOtDwYHWiStizrdRHVA/v0TLLmT97HxSSOeUGlbycyMi7PjKtRnCqmLJOZDmhw
I0OQsiJC+/lQST60krBmTAL9FzuNayfNVTEAlsGiifXrnHQTjtKBjo1F245/Q6FD
MyD80oZ6zoCVvd+jlV2CD44wurnvihZIU6UQXxXscniF5hvFVEdBZoR7C8YoFb/4
VCMOX+Et4SfA3l9HwldAEj9HndGxtYXthrmmOt6TUiK6hBAPdrTCnKDmmMruraDS
pGzKCkVWg84FV5fGekt4MYJWAsA3pX0Bbp/9xnXAGJpEPS+bMSp6Fb+paZ6oFd49
EJtmkI4pWNHbGYQSYcHQAisuve5uLshcaz5XOc20j3JaC4N6kQ8rjbnRjhRjYkle
jO0e1MnkWCJohTw2C2s4AR1iYir+6Do4I9a7fAy7XdwhCaME9rqnWSFu4YqY60TV
8v/cuYe143zIhwiQg8I3nxNEKK24qSFucCpiGnfSU+ZxP7IAnN0TUl5KW8FitFOJ
rLuUlpSsC+sOBo17tepcuZrYNzg33d5h9Y5swRaQsYCaMf0HaiovijJ2D+qU9Dbc
yS9aoDWmh3Uzh16W+FeyGszjpgF2WUhtl25Z87Nyi2eCLsd1ndRzRNx1EUy+M2iv
OLGzktQ7aQ47rYlSekhUclsACw6II3hsfBiyQvp01LtGEe54YjIcMM33LQ2yEl2l
sZCwcM3aXcy851TqPNvcTRg8OHeW+4soGmYLAIIqs4CJ4oss2ei9RTMDflCML0av
AZOz+H28aOggZsiVheclkV0gC3dMeH9SHpD7OxgKnWWIBFmOHO18mHan5zS4LEaw
vvhJkQC44WR+aoiZtfWicFGKD7ylBuGalg6V7lrij6viYd0atCfgJM/6ZhxtO8e2
SjJMPTqf/W6Wvgl07yBHZEqTkoT3yo0/sUXlcJ5yIhAOmE5ONu4RkoXvH3cYP1so
f0kXIfeCOderYK3f9wMU3ND8w7EZzbTe/gPz9Sis/4lKsJ2OND+0ZA4711e5S44T
dNSxeeaIFeMJFMYKSOzCbCo3PatyfzQCIHwvvDWjv69manSvG49v0wEnMpEwNbMJ
hFNAFaES+G0ENDdFHYON/RTrlePVAuFUpV4WmMrC5UWDoG9bP17s2ITotbvgk3wG
ZpeRVFVU4GiRJw/m/H7GUXZsl4maCm8N4Xi74FKXlMPC3vbnSjYu1OM1/L/8MI+E
R8URJxS2+/F6E4jmgEADmWREVQVP2RNFO3xmMBPYDdl2NK+ADJATMobphC09StQ7
LpkY6/3P+WQvax2P9RKefuuA6fIe6/o8WOaoASLheOitzqgICa6WnuGd7I0kqjNq
sCBkZGHLOtJpxHXloVcMKztAIaEFGnOUeGZYQw1eUpscqY9c/XB0uWiyx6JBNnID
4doyn3RYihW0ji+hJCSvaUS2UEUCAdMpigjWMHYrfb8+Zbfd+LCQUCFPmQ7Y9YwD
DoIbDnsn/iTavbfepVL0yf7xEIunOA1vWIzcNMQ6bu/a06+aAAinhpZhqLrz9bcz
p0hBwVo4IB9a7X6kaD6bqzb2I64npdUr+gW5yaUhZ5iKpCpaMOIuREUFOaD2RV71
slMiKo8Axdj0hTzYsyY3t0NeyxbG4+M6eAB4avz+8sDfD+JnsZqzG4alK45wnQG2
zEW9zG3FMrnifL1c6rDYuM8bFmCYfQn2dX63FClgcQv7Mw+iBFLMto2+w0oMkWhj
60eLRFlJZDDNxCM1DdxE+tRP9Ju/svCuJQAWrTzP5BfhCOL4ojXix52WRNnpYohy
sPmamrD1VmY937k2WIQ9Xi3G5WEEWJqH2Q+jPFehLnnSF+cVxQB8J5GC7j+pO/sv
uFojUCgIDq78Ap7nqCNUGbb8gWKJFJN2TtqvA/rrZadPPktdMNtBDHX1hS5ZI+1N
b5X7gtYPNZvJacIYoS9gLxQv9U6LficaXtGvJXrlr32hcXk+jAw79ViGzmIU3TsY
ltp1UKgoo8deIs+m9qzkKT5votmfUdlcgdNuqpRVXe4Qv5TljI9HjC3P92epdlLr
8BoT7gfy4g==
